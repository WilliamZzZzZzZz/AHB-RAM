`ifndef AHBRAM_SMOKE_TEST_SV
`define AHBRAM_SMOKE_TEST_SV

class ahbram_smoke_test extends ahbram_base_test;

    `uvm_component_utils(ahbram_smoke_test)

    function new(string name = "ahbram_smoke_test", uvm_componemnt parent);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
    endfunction

    task run_phase(uvm_phase phase);
        ahbram_smoke_virtual_sequence seq = ahbram_smoke_virtual_sequence::type_id::create("seq");
        super.run_phase(phase);

        phase.raise_objection(this);
        seq.start(env.virt_sqr);
        phase.drop_objection(this);
        
    endtask


endclass

`endif 