`ifndef AHBRAM_PKG_SV
`define AHBRAM_PKG_SV

package my_uvm_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import ahb_pkg::*;

    `include "ahbram_configuration.sv"
    `include "ahbram_env.sv"
    `include "ahbram_scoreboard.sv"
    `include "ahbram_subscriber.sv"
    `include "ahbram_virtual_sequencer.sv"

    `include "ahbram_element_sequences.svh"
    `include "ahbram_sequence_lib.svh"
    `include "ahbram_tests.svh"

endpackage

`endif 