`ifndef AHBRAM_TESTS_SV
`define AHBRAM_TSETS_SV

`include "ahbram_base_test.sv"
`include "ahbram_smoke_test.sv"

`endif 