`ifndef AHBRAM_IF_SV
`define AHBRAM_IF_SV

interface ahbram_if;

endinterface

`endif 