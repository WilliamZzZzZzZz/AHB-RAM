`ifndef AHBRAM_SEQUENCE_LIB_SVH
`define AHBRAM_SEQUENCE_LIB_SVH

`include "ahbram_element_sequences.svh"
`include "ahbram_base_virtual_sequence.sv"
`include "ahbram_smoke_virtual_sequence.sv"

`endif 