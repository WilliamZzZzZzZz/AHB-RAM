`ifndef AHB_MASTER_AGENT_SV
`define AHB_MASTER_AGENT_SV

class ahb_master_agent extends uvm_agent;

    ahb_agent_configuration cfg;

    ahb_master_driver

endclass

`endif 