`ifndef AHBRAM_ELEMENT_SEQUENCES_SV
`define AHBRAM_ELEMENT_SEQUENCES_SV

`include "ahbram_base_element_sequence.sv"
`include "ahbram_single_read_sequence.sv"
`include "ahbram_single_write_sequence.sv"

`endif 