`ifndef AHB_IF_SV
`define AHB_IF_SV

interface ahb_if;

endinterface

`endif 